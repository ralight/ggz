<div id="acknowledgements">
	<div class="note" style="float:left;">
		&copy; 2005 <a href="http://www.ggzgamingzone.org/">GGZ Gaming Zone</a>
	</div>
	<div class="note" style="float:right;">
		Design baserad på Steel-n-Leather &copy; 2004 av
		<a href="mailto:brian.allbee@gmail.com" title="Comment on this design if you wish!">Brian D. Allbee</a>
	</div>
	<div class="note" style="float:left;">
	<?php
		Locale::availablelanguages();
	?>
	</div>
</div>
