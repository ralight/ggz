	<div class="menubar">
		<div class="menu">
			<a href="/" class="menuitem" title="Startsida">Start</a>
		</div>
		<div class="menu">
			<a href="/db/" class="menuitem" title="Spelstatistik och rank">Databas</a>
			<div class="menu">
				<a href="/db/" class="menuitem">Överblick</a>
				<a href="/db/games/" class="menuitem">Spel</a>
				<a href="/db/matches/" class="menuitem">Matcher</a>
				<a href="/db/tournaments/" class="menuitem">Turneringar</a>
				<a href="/db/players/" class="menuitem">Spelare</a>
				<a href="/db/teams/" class="menuitem">Teams/Klaner</a>
			</div>
		</div>
		<div class="menu">
			<a href="/games/" class="menuitem" title="Lite online-kul">Spela!</a>
			<div class="menu">
				<a href="/games/" class="menuitem">GGZ-spel</a>
				<a href="/webgames/" class="menuitem">Web-spel</a>
			</div>
		</div>
		<div class="menu">
			<a href="/active/hotstuff/" class="menuitem" title="Användarbidrag">Organisera!</a>
			<div class="menu">
				<a href="/active/hotstuff/" class="menuitem">Spel-innehåll</a>
				<a href="/active/tournaments/" class="menuitem">Turneringar</a>
				<a href="/active/teams/" class="menuitem">Teams/Klaner</a>
			</div>
		</div>
		<div class="menu">
			<a href="/forums/" class="menuitem" title="Forum">Forum</a>
			<div class="menu">
				<a href="/forums/" class="menuitem">Kommunity-forum</a>
				<a href="/blogs/" class="menuitem">Individuella bloggar</a>
				<a href="/articles/" class="menuitem">Artiklar</a>
			</div>
		</div>
		<div class="menu">
			<a href="/contact/" class="menuitem" title="Om GGZ-Kommunity">Om</a>
			<div class="menu">
				<a href="/contact/" class="menuitem">Kontakt</a>
			</div>
		</div>
	</div>
