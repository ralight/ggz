	<div style="float:left">
	<img src="<?php Config::theme("pagelogo.png"); ?>" alt="Community logo">
	</div>
	<div style="margin-top: 8px">
	<h1>GGZ Kommunity</h1>
	<h2>Spelportalen baserad på GGZ Gaming Zone</h2>
	</div>
