<div id="main">
	<h1>
		<span class="itemleader">:: </span>
		Programming for GGZ in Ruby
		<span class="itemleader"> :: </span>
		<a name="ruby"></a>
	</h1>
	<div class="text">
		<div style="float:right">
		<img src="images/ruby.png" alt="Ruby logo">
		</div>
		While development in C, C++ and Python has been possible for a long time
		already, some progress has recently been experienced with reviving the old
		Ruby bindings of GGZ.
		For the time being, a simple GGZdMod wrapper exists, which has been used
		to implement an alternative Tic-Tac-Toe server, sharing the AI routines
		with the original one. Read about it in our article:
		<a href="/articles/ruby/" title="GGZ and Ruby">GGZ and Ruby</a>.
	</div>

	<h1>
		<span class="itemleader">:: </span>
		Extending the Community platform
		<span class="itemleader"> :: </span>
		<a name="extending"></a>
	</h1>
	<div class="text">
		The GGZ Community portal is being extended so it can be used more easily
		by other projects as well. This includes custom stylesheets, internationalization
		and a template and configuration system.
		If anyone wants to help with the translation, the current message catalog is
		as usually available
		<a href="http://dev.ggzgamingzone.org/i18n/" title="GGZ Internationalization">on our i18n page</a>, and takes up about 100 strings out of 2200 which GGZ has in total.
	</div>

	<h1>
		<span class="itemleader">:: </span>
		GGZ 0.0.11 and Packaging article
		<span class="itemleader"> :: </span>
		<a name="0011"></a>
	</h1>
	<div class="text">
		<div style="float:left">
		<img src="images/packagesarticle.png" alt="GGZ package overview">
		</div>
		You can now <a href="http://www.ggzgamingzone.org/">download</a>
		GGZ 0.0.11 from the project site, and if you're a packager,
		do not miss our new article:
		<a href="/articles/packaging/" title="GGZ packaging">GGZ packaging</a>.
	</div>

	<h1>
		<span class="itemleader">:: </span>
		Server move and updates
		<span class="itemleader"> :: </span>
		<a name="servermove"></a>
	</h1>
	<div class="text">
		The GGZ Community has moved off the project server and to another
		dedicated server located in France. We're using the chance on upgrading
		it to the current CVS version. This brings along with it longitude/latitude
		configuration in the personal settings (for the world map), a karma
		system, and preparations for the upcoming GGZ release's savegames.
	</div>

	<h1>
		<span class="itemleader">:: </span>
		GGZ Gaming Zone 0.0.10 released
		<span class="itemleader"> :: </span>
		<a name="0010"></a>
	</h1>
	<div class="text">
		Version 0.0.10 of the GGZ project had been released last night (24.01.2005).
		Information about it can be found at the release announcement
		<a href="http://www.ggzgamingzone.org/releases/0.0.10/release.php">page</a>.
		A couple of new games have been installed and are now moving into the
		database of already played games
		(<a href="/db/games/?lookup=Hnefatafl" title="Hnefatafl">Hnefatafl</a>,
		<a href="/db/games/?lookup=Checkers" title="Dame">Checkers</a>,
		<a href="/db/games/?lookup=Krosswater" title="Krosswater">Krosswater</a>).
		Do not forget to add your blogs to the
		<a href="/blogs/" title="Planet GGZ Community">Blog collection</a>.
		Have fun :)
	</div>

	<h1>
		<span class="itemleader">:: </span>
		Jubileum: 5 år av GGZ Gaming Zone!
		<span class="itemleader"> :: </span>
		<a name="5years"></a>
	</h1>
	<div class="text">
		<div style="float:right">
		<img src="images/grubbyparty.png" alt="Grubby bjuder in dej!">
		</div>
		Det är otroligt - projektet blev 5 år gammalt idag!
		Ta en titt på den speciellt tillägnade
		<a href="/5years/" title="GGZs femte födelsedag">födelsedagssidan</a>.
	</div>

	<h1>
		<span class="itemleader">:: </span>
		Ny GGZ-Kommunityportal
		<span class="itemleader"> ::</span>
		<a name="newportal"></a>
	</h1>
	<div class="text">
		Ersätter de gamla <a href="http://www.ggzgamingzone.org/backend/web/" title="">Ranking</a>
		-sidorna, och siktar på mycket mer:
		Statistik om allt spelrelaterat på GGZ, användarinsända nivåer och teman, forum och
		bloggar, spelrecensioner, organiserade turneringar, och små underhållande webspel.
		GGZ-servrar kan använda "ggz-community" paketet för att göra egna portaler.
	</div>

</div>
