<?php include("top.inc"); ?>

<div id="main">
	<h1>
		<span class="itemleader">:: </span>
		Om GGZ-Kommunityportalen
		<span class="itemleader"> :: </span>
		<a name="about"></a>
	</h1>
	<div class="text">
		<div>
		Firandes sin femte födelsedag, har
		<a href="http://www.ggzgamingzone.org/">GGZ Gaming Zone</a>
		-projektet invigt GGZ Kommunity, en portal tillägnad
		spelare (och blivande spelare) av GGZ-spel.
		</div>
	</div>

	<h1>
		<span class="itemleader">:: </span>
		Kontakta oss
		<span class="itemleader"> ::</span>
		<a name="contact"></a>
	</h1>
	<div class="text">
		Du kan skicka oss epost när helst du önskar, förutom spam
		förståss :)
		<br>
		Addresen är:
		<a href="mailto:info@ggzcommunity.org">info@ggzcommunity.org</a>
		<br><br>
		För frågor angående utvecklandet av GGZ, ta en titt på projektets
		<a href="https://mail.ggzgamingzone.org/">mejllistor</a>.
	</div>

</div>

<?php include("bottom.inc"); ?>
